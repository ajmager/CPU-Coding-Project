//datapath.v
module datapath (clr, );