library verilog;
use verilog.vl_types.all;
entity datapath is
    port(
        clk             : in     vl_logic;
        clr             : in     vl_logic;
        r0_in           : in     vl_logic;
        r1_in           : in     vl_logic;
        r2_in           : in     vl_logic;
        r3_in           : in     vl_logic;
        r4_in           : in     vl_logic;
        r5_in           : in     vl_logic;
        r6_in           : in     vl_logic;
        r7_in           : in     vl_logic;
        r8_in           : in     vl_logic;
        r9_in           : in     vl_logic;
        r10_in          : in     vl_logic;
        r11_in          : in     vl_logic;
        r12_in          : in     vl_logic;
        r13_in          : in     vl_logic;
        r14_in          : in     vl_logic;
        r15_in          : in     vl_logic;
        PC_in           : in     vl_logic;
        Inc_PC          : in     vl_logic;
        IR_in           : in     vl_logic;
        Y_in            : in     vl_logic;
        Z_in            : in     vl_logic;
        HI_in           : in     vl_logic;
        LO_in           : in     vl_logic;
        MAR_in          : in     vl_logic;
        MDR_in          : in     vl_logic;
        read            : in     vl_logic;
        inPort_in       : in     vl_logic;
        r0out           : in     vl_logic;
        r1out           : in     vl_logic;
        r2out           : in     vl_logic;
        r3out           : in     vl_logic;
        r4out           : in     vl_logic;
        r5out           : in     vl_logic;
        r6out           : in     vl_logic;
        r7out           : in     vl_logic;
        r8out           : in     vl_logic;
        r9out           : in     vl_logic;
        r10out          : in     vl_logic;
        r11out          : in     vl_logic;
        r12out          : in     vl_logic;
        r13out          : in     vl_logic;
        r14out          : in     vl_logic;
        r15out          : in     vl_logic;
        PCout           : in     vl_logic;
        ZLOWout         : in     vl_logic;
        ZHIout          : in     vl_logic;
        LOout           : in     vl_logic;
        HIout           : in     vl_logic;
        MDRout          : in     vl_logic;
        inPortout       : in     vl_logic;
        Cout            : in     vl_logic;
        ALU_select      : in     vl_logic_vector(3 downto 0);
        MdataIn         : in     vl_logic_vector(31 downto 0);
        ALU_out         : out    vl_logic_vector(63 downto 0)
    );
end datapath;
