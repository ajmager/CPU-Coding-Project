library verilog;
use verilog.vl_types.all;
entity \bus\ is
    port(
        r0_out          : in     vl_logic_vector(31 downto 0);
        r1_out          : in     vl_logic_vector(31 downto 0);
        r2_out          : in     vl_logic_vector(31 downto 0);
        r3_out          : in     vl_logic_vector(31 downto 0);
        r4_out          : in     vl_logic_vector(31 downto 0);
        r5_out          : in     vl_logic_vector(31 downto 0);
        r6_out          : in     vl_logic_vector(31 downto 0);
        r7_out          : in     vl_logic_vector(31 downto 0);
        r8_out          : in     vl_logic_vector(31 downto 0);
        r9_out          : in     vl_logic_vector(31 downto 0);
        r10_out         : in     vl_logic_vector(31 downto 0);
        r11_out         : in     vl_logic_vector(31 downto 0);
        r12_out         : in     vl_logic_vector(31 downto 0);
        r13_out         : in     vl_logic_vector(31 downto 0);
        r14_out         : in     vl_logic_vector(31 downto 0);
        r15_out         : in     vl_logic_vector(31 downto 0);
        HI_out          : in     vl_logic_vector(31 downto 0);
        LO_out          : in     vl_logic_vector(31 downto 0);
        ZHI_out         : in     vl_logic_vector(31 downto 0);
        ZLOW_out        : in     vl_logic_vector(31 downto 0);
        PC_out          : in     vl_logic_vector(31 downto 0);
        MDR_out         : in     vl_logic_vector(31 downto 0);
        inPort_out      : in     vl_logic_vector(31 downto 0);
        C_sign_extended : in     vl_logic_vector(31 downto 0);
        r0out           : in     vl_logic;
        r1out           : in     vl_logic;
        r2out           : in     vl_logic;
        r3out           : in     vl_logic;
        r4out           : in     vl_logic;
        r5out           : in     vl_logic;
        r6out           : in     vl_logic;
        r7out           : in     vl_logic;
        r8out           : in     vl_logic;
        r9out           : in     vl_logic;
        r10out          : in     vl_logic;
        r11out          : in     vl_logic;
        r12out          : in     vl_logic;
        r13out          : in     vl_logic;
        r14out          : in     vl_logic;
        r15out          : in     vl_logic;
        HIout           : in     vl_logic;
        LOout           : in     vl_logic;
        ZHIout          : in     vl_logic;
        ZLOWout         : in     vl_logic;
        PCout           : in     vl_logic;
        MDRout          : in     vl_logic;
        inPortout       : in     vl_logic;
        Cout            : in     vl_logic;
        BUS_data        : out    vl_logic_vector(31 downto 0);
        clk             : in     vl_logic
    );
end \bus\;
